//****** set a PARAMETER_DATA_MODE setting to "D" / DATA_MODE = "R"
//****** add a TEMP_DOXY_ADJUSTED value in an to a "R" variable *****

netcdf BR1900722_002 {
dimensions:
	DATE_TIME = 14 ;
	STRING2 = 2 ;
	STRING4 = 4 ;
	STRING8 = 8 ;
	STRING16 = 16 ;
	STRING32 = 32 ;
	STRING64 = 64 ;
	STRING256 = 256 ;
	N_PROF = 1 ;
	N_PARAM = 4 ;
	N_LEVELS = 71 ;
	N_CALIB = 1 ;
	N_HISTORY = UNLIMITED ; // (1 currently)
variables:
	char DATA_TYPE(STRING32) ;
		DATA_TYPE:long_name = "Data type" ;
		DATA_TYPE:conventions = "Argo reference table 1" ;
		DATA_TYPE:_FillValue = " " ;
	char FORMAT_VERSION(STRING4) ;
		FORMAT_VERSION:long_name = "File format version" ;
		FORMAT_VERSION:_FillValue = " " ;
	char HANDBOOK_VERSION(STRING4) ;
		HANDBOOK_VERSION:long_name = "Data handbook version" ;
		HANDBOOK_VERSION:_FillValue = " " ;
	char REFERENCE_DATE_TIME(DATE_TIME) ;
		REFERENCE_DATE_TIME:long_name = "Date of reference for Julian days" ;
		REFERENCE_DATE_TIME:conventions = "YYYYMMDDHHMISS" ;
		REFERENCE_DATE_TIME:_FillValue = " " ;
	char PLATFORM_NUMBER(N_PROF, STRING8) ;
		PLATFORM_NUMBER:long_name = "Float unique identifier" ;
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII" ;
		PLATFORM_NUMBER:_FillValue = " " ;
	char PROJECT_NAME(N_PROF, STRING64) ;
		PROJECT_NAME:long_name = "Name of the project" ;
		PROJECT_NAME:_FillValue = " " ;
	char PI_NAME(N_PROF, STRING64) ;
		PI_NAME:long_name = "Name of the principal investigator" ;
		PI_NAME:_FillValue = " " ;
	char STATION_PARAMETERS(N_PROF, N_PARAM, STRING64) ;
		STATION_PARAMETERS:long_name = "List of available parameters for the station" ;
		STATION_PARAMETERS:conventions = "Argo reference table 3" ;
		STATION_PARAMETERS:_FillValue = " " ;
	int CYCLE_NUMBER(N_PROF) ;
		CYCLE_NUMBER:long_name = "Float cycle number" ;
		CYCLE_NUMBER:conventions = "0...N, 0 : launch cycle (if exists), 1 : first complete cycle" ;
		CYCLE_NUMBER:_FillValue = 99999 ;
	char DIRECTION(N_PROF) ;
		DIRECTION:long_name = "Direction of the station profiles" ;
		DIRECTION:conventions = "A: ascending profiles, D: descending profiles" ;
		DIRECTION:_FillValue = " " ;
	char DATA_CENTRE(N_PROF, STRING2) ;
		DATA_CENTRE:long_name = "Data centre in charge of float data processing" ;
		DATA_CENTRE:conventions = "Argo reference table 4" ;
		DATA_CENTRE:_FillValue = " " ;
	char DATE_CREATION(DATE_TIME) ;
		DATE_CREATION:long_name = "Date of file creation" ;
		DATE_CREATION:conventions = "YYYYMMDDHHMISS" ;
		DATE_CREATION:_FillValue = " " ;
	char DATE_UPDATE(DATE_TIME) ;
		DATE_UPDATE:long_name = "Date of update of this file" ;
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS" ;
		DATE_UPDATE:_FillValue = " " ;
	char DC_REFERENCE(N_PROF, STRING32) ;
		DC_REFERENCE:long_name = "Station unique identifier in data centre" ;
		DC_REFERENCE:conventions = "Data centre convention" ;
		DC_REFERENCE:_FillValue = " " ;
	char DATA_STATE_INDICATOR(N_PROF, STRING4) ;
		DATA_STATE_INDICATOR:long_name = "Degree of processing the data have passed through" ;
		DATA_STATE_INDICATOR:conventions = "Argo reference table 6" ;
		DATA_STATE_INDICATOR:_FillValue = " " ;
	char DATA_MODE(N_PROF) ;
		DATA_MODE:long_name = "Delayed mode or real time data" ;
		DATA_MODE:conventions = "R : real time; D : delayed mode; A : real time with adjustment" ;
		DATA_MODE:_FillValue = " " ;
	char PARAMETER_DATA_MODE(N_PROF, N_PARAM) ;
		PARAMETER_DATA_MODE:long_name = "Delayed mode or real time data" ;
		PARAMETER_DATA_MODE:conventions = "R : real time; D : delayed mode; A : real time with adjustment" ;
		PARAMETER_DATA_MODE:_FillValue = " " ;
	char PLATFORM_TYPE(N_PROF, STRING32) ;
		PLATFORM_TYPE:long_name = "Type of float" ;
		PLATFORM_TYPE:conventions = "Argo reference table 23" ;
		PLATFORM_TYPE:_FillValue = " " ;
	char FLOAT_SERIAL_NO(N_PROF, STRING32) ;
		FLOAT_SERIAL_NO:long_name = "Serial number of the float" ;
		FLOAT_SERIAL_NO:_FillValue = " " ;
	char FIRMWARE_VERSION(N_PROF, STRING32) ;
		FIRMWARE_VERSION:long_name = "Instrument firmware version" ;
		FIRMWARE_VERSION:_FillValue = " " ;
	char WMO_INST_TYPE(N_PROF, STRING4) ;
		WMO_INST_TYPE:long_name = "Coded instrument type" ;
		WMO_INST_TYPE:conventions = "Argo reference table 8" ;
		WMO_INST_TYPE:_FillValue = " " ;
	double JULD(N_PROF) ;
		JULD:long_name = "Julian day (UTC) of the station relative to REFERENCE_DATE_TIME" ;
		JULD:standard_name = "time" ;
		JULD:units = "days since 1950-01-01 00:00:00 UTC" ;
		JULD:conventions = "Relative julian days with decimal part (as parts of day)" ;
		JULD:resolution = 1.e-08 ;
		JULD:_FillValue = 999999. ;
		JULD:axis = "T" ;
	char JULD_QC(N_PROF) ;
		JULD_QC:long_name = "Quality on date and time" ;
		JULD_QC:conventions = "Argo reference table 2" ;
		JULD_QC:_FillValue = " " ;
	double JULD_LOCATION(N_PROF) ;
		JULD_LOCATION:long_name = "Julian day (UTC) of the location relative to REFERENCE_DATE_TIME" ;
		JULD_LOCATION:units = "days since 1950-01-01 00:00:00 UTC" ;
		JULD_LOCATION:conventions = "Relative julian days with decimal part (as parts of day)" ;
		JULD_LOCATION:resolution = 1.e-08 ;
		JULD_LOCATION:_FillValue = 999999. ;
	double LATITUDE(N_PROF) ;
		LATITUDE:long_name = "Latitude of the station, best estimate" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degree_north" ;
		LATITUDE:_FillValue = 99999. ;
		LATITUDE:valid_min = -90. ;
		LATITUDE:valid_max = 90. ;
		LATITUDE:axis = "Y" ;
	double LONGITUDE(N_PROF) ;
		LONGITUDE:long_name = "Longitude of the station, best estimate" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degree_east" ;
		LONGITUDE:_FillValue = 99999. ;
		LONGITUDE:valid_min = -180. ;
		LONGITUDE:valid_max = 180. ;
		LONGITUDE:axis = "X" ;
	char POSITION_QC(N_PROF) ;
		POSITION_QC:long_name = "Quality on position (latitude and longitude)" ;
		POSITION_QC:conventions = "Argo reference table 2" ;
		POSITION_QC:_FillValue = " " ;
	char POSITIONING_SYSTEM(N_PROF, STRING8) ;
		POSITIONING_SYSTEM:long_name = "Positioning system" ;
		POSITIONING_SYSTEM:_FillValue = " " ;
	char VERTICAL_SAMPLING_SCHEME(N_PROF, STRING256) ;
		VERTICAL_SAMPLING_SCHEME:long_name = "Vertical sampling scheme" ;
		VERTICAL_SAMPLING_SCHEME:conventions = "Argo reference table 16" ;
		VERTICAL_SAMPLING_SCHEME:_FillValue = " " ;
	int CONFIG_MISSION_NUMBER(N_PROF) ;
		CONFIG_MISSION_NUMBER:long_name = "Unique number denoting the missions performed by the float" ;
		CONFIG_MISSION_NUMBER:conventions = "1...N, 1 : first complete mission" ;
		CONFIG_MISSION_NUMBER:_FillValue = 99999 ;
	char PROFILE_TEMP_DOXY_QC(N_PROF) ;
		PROFILE_TEMP_DOXY_QC:long_name = "Global quality flag of TEMP_DOXY profile" ;
		PROFILE_TEMP_DOXY_QC:conventions = "Argo reference table 2a" ;
		PROFILE_TEMP_DOXY_QC:_FillValue = " " ;
	char PROFILE_BPHASE_DOXY_QC(N_PROF) ;
		PROFILE_BPHASE_DOXY_QC:long_name = "Global quality flag of BPHASE_DOXY profile" ;
		PROFILE_BPHASE_DOXY_QC:conventions = "Argo reference table 2a" ;
		PROFILE_BPHASE_DOXY_QC:_FillValue = " " ;
	char PROFILE_DOXY_QC(N_PROF) ;
		PROFILE_DOXY_QC:long_name = "Global quality flag of DOXY profile" ;
		PROFILE_DOXY_QC:conventions = "Argo reference table 2a" ;
		PROFILE_DOXY_QC:_FillValue = " " ;
	float PRES(N_PROF, N_LEVELS) ;
		PRES:long_name = "Sea water pressure, equals 0 at sea-level" ;
		PRES:standard_name = "sea_water_pressure" ;
		PRES:units = "decibar" ;
		PRES:valid_min = 0.f ;
		PRES:valid_max = 12000.f ;
		PRES:resolution = 0.1f ;
		PRES:C_format = "%7.1f" ;
		PRES:FORTRAN_format = "F7.1f" ;
		PRES:_FillValue = 99999.f ;
		PRES:axis = "Z" ;
	float TEMP_DOXY(N_PROF, N_LEVELS) ;
		TEMP_DOXY:long_name = "Sea temperature from oxygen sensor ITS-90 scale" ;
		TEMP_DOXY:standard_name = "temperature_of_sensor_for_oxygen_in_sea_water" ;
		TEMP_DOXY:units = "degree_Celsius" ;
		TEMP_DOXY:valid_min = -2.f ;
		TEMP_DOXY:valid_max = 40.f ;
		TEMP_DOXY:resolution = 0.001f ;
		TEMP_DOXY:C_format = "%9.3f" ;
		TEMP_DOXY:FORTRAN_format = "F9.3f" ;
		TEMP_DOXY:_FillValue = 99999.f ;
	char TEMP_DOXY_QC(N_PROF, N_LEVELS) ;
		TEMP_DOXY_QC:long_name = "quality flag" ;
		TEMP_DOXY_QC:conventions = "Argo reference table 2" ;
		TEMP_DOXY_QC:_FillValue = " " ;
	float TEMP_DOXY_ADJUSTED(N_PROF, N_LEVELS) ;
		TEMP_DOXY_ADJUSTED:long_name = "Sea temperature from oxygen sensor ITS-90 scale" ;
		TEMP_DOXY_ADJUSTED:standard_name = "temperature_of_sensor_for_oxygen_in_sea_water" ;
		TEMP_DOXY_ADJUSTED:units = "degree_Celsius" ;
		TEMP_DOXY_ADJUSTED:valid_min = -2.f ;
		TEMP_DOXY_ADJUSTED:valid_max = 40.f ;
		TEMP_DOXY_ADJUSTED:resolution = 0.001f ;
		TEMP_DOXY_ADJUSTED:C_format = "%9.3f" ;
		TEMP_DOXY_ADJUSTED:FORTRAN_format = "F9.3f" ;
		TEMP_DOXY_ADJUSTED:_FillValue = 99999.f ;
	char TEMP_DOXY_ADJUSTED_QC(N_PROF, N_LEVELS) ;
		TEMP_DOXY_ADJUSTED_QC:long_name = "quality flag" ;
		TEMP_DOXY_ADJUSTED_QC:conventions = "Argo reference table 2" ;
		TEMP_DOXY_ADJUSTED_QC:_FillValue = " " ;
	float TEMP_DOXY_ADJUSTED_ERROR(N_PROF, N_LEVELS) ;
		TEMP_DOXY_ADJUSTED_ERROR:long_name = "Contains the error on the adjusted values as determined by the delayed mode QC process" ;
		TEMP_DOXY_ADJUSTED_ERROR:units = "degree_Celsius" ;
		TEMP_DOXY_ADJUSTED_ERROR:resolution = 0.001f ;
		TEMP_DOXY_ADJUSTED_ERROR:C_format = "%9.3f" ;
		TEMP_DOXY_ADJUSTED_ERROR:FORTRAN_format = "F9.3f" ;
		TEMP_DOXY_ADJUSTED_ERROR:_FillValue = 99999.f ;
	float BPHASE_DOXY(N_PROF, N_LEVELS) ;
		BPHASE_DOXY:long_name = "Uncalibrated phase shift reported by oxygen sensor" ;
		BPHASE_DOXY:units = "degree" ;
		BPHASE_DOXY:valid_min = 10.f ;
		BPHASE_DOXY:valid_max = 70.f ;
		BPHASE_DOXY:resolution = 0.01f ;
		BPHASE_DOXY:C_format = "%8.2f" ;
		BPHASE_DOXY:FORTRAN_format = "F8.2f" ;
		BPHASE_DOXY:_FillValue = 99999.f ;
	char BPHASE_DOXY_QC(N_PROF, N_LEVELS) ;
		BPHASE_DOXY_QC:long_name = "quality flag" ;
		BPHASE_DOXY_QC:conventions = "Argo reference table 2" ;
		BPHASE_DOXY_QC:_FillValue = " " ;
	float BPHASE_DOXY_ADJUSTED(N_PROF, N_LEVELS) ;
		BPHASE_DOXY_ADJUSTED:long_name = "Uncalibrated phase shift reported by oxygen sensor" ;
		BPHASE_DOXY_ADJUSTED:units = "degree" ;
		BPHASE_DOXY_ADJUSTED:valid_min = 10.f ;
		BPHASE_DOXY_ADJUSTED:valid_max = 70.f ;
		BPHASE_DOXY_ADJUSTED:resolution = 0.01f ;
		BPHASE_DOXY_ADJUSTED:C_format = "%8.2f" ;
		BPHASE_DOXY_ADJUSTED:FORTRAN_format = "F8.2f" ;
		BPHASE_DOXY_ADJUSTED:_FillValue = 99999.f ;
	char BPHASE_DOXY_ADJUSTED_QC(N_PROF, N_LEVELS) ;
		BPHASE_DOXY_ADJUSTED_QC:long_name = "quality flag" ;
		BPHASE_DOXY_ADJUSTED_QC:conventions = "Argo reference table 2" ;
		BPHASE_DOXY_ADJUSTED_QC:_FillValue = " " ;
	float BPHASE_DOXY_ADJUSTED_ERROR(N_PROF, N_LEVELS) ;
		BPHASE_DOXY_ADJUSTED_ERROR:long_name = "Contains the error on the adjusted values as determined by the delayed mode QC process" ;
		BPHASE_DOXY_ADJUSTED_ERROR:units = "degree" ;
		BPHASE_DOXY_ADJUSTED_ERROR:resolution = 0.01f ;
		BPHASE_DOXY_ADJUSTED_ERROR:C_format = "%8.2f" ;
		BPHASE_DOXY_ADJUSTED_ERROR:FORTRAN_format = "F8.2f" ;
		BPHASE_DOXY_ADJUSTED_ERROR:_FillValue = 99999.f ;
	float DOXY(N_PROF, N_LEVELS) ;
		DOXY:long_name = "Dissolved oxygen" ;
		DOXY:standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water" ;
		DOXY:units = "micromole/kg" ;
		DOXY:valid_min = 0.f ;
		DOXY:valid_max = 600.f ;
		DOXY:resolution = 0.001f ;
		DOXY:C_format = "%9.3f" ;
		DOXY:FORTRAN_format = "F9.3f" ;
		DOXY:_FillValue = 99999.f ;
	char DOXY_QC(N_PROF, N_LEVELS) ;
		DOXY_QC:long_name = "quality flag" ;
		DOXY_QC:conventions = "Argo reference table 2" ;
		DOXY_QC:_FillValue = " " ;
	float DOXY_ADJUSTED(N_PROF, N_LEVELS) ;
		DOXY_ADJUSTED:long_name = "Dissolved oxygen" ;
		DOXY_ADJUSTED:standard_name = "moles_of_oxygen_per_unit_mass_in_sea_water" ;
		DOXY_ADJUSTED:units = "micromole/kg" ;
		DOXY_ADJUSTED:valid_min = 0.f ;
		DOXY_ADJUSTED:valid_max = 600.f ;
		DOXY_ADJUSTED:resolution = 0.001f ;
		DOXY_ADJUSTED:C_format = "%9.3f" ;
		DOXY_ADJUSTED:FORTRAN_format = "F9.3f" ;
		DOXY_ADJUSTED:_FillValue = 99999.f ;
	char DOXY_ADJUSTED_QC(N_PROF, N_LEVELS) ;
		DOXY_ADJUSTED_QC:long_name = "quality flag" ;
		DOXY_ADJUSTED_QC:conventions = "Argo reference table 2" ;
		DOXY_ADJUSTED_QC:_FillValue = " " ;
	float DOXY_ADJUSTED_ERROR(N_PROF, N_LEVELS) ;
		DOXY_ADJUSTED_ERROR:long_name = "Contains the error on the adjusted values as determined by the delayed mode QC process" ;
		DOXY_ADJUSTED_ERROR:units = "micromole/kg" ;
		DOXY_ADJUSTED_ERROR:resolution = 0.001f ;
		DOXY_ADJUSTED_ERROR:C_format = "%9.3f" ;
		DOXY_ADJUSTED_ERROR:FORTRAN_format = "F9.3f" ;
		DOXY_ADJUSTED_ERROR:_FillValue = 99999.f ;
	char PARAMETER(N_PROF, N_CALIB, N_PARAM, STRING64) ;
		PARAMETER:long_name = "List of parameters with calibration information" ;
		PARAMETER:conventions = "Argo reference table 3" ;
		PARAMETER:_FillValue = " " ;
	char SCIENTIFIC_CALIB_EQUATION(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_EQUATION:long_name = "Calibration equation for this parameter" ;
		SCIENTIFIC_CALIB_EQUATION:_FillValue = " " ;
	char SCIENTIFIC_CALIB_COEFFICIENT(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_COEFFICIENT:long_name = "Calibration coefficients for this equation" ;
		SCIENTIFIC_CALIB_COEFFICIENT:_FillValue = " " ;
	char SCIENTIFIC_CALIB_COMMENT(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_COMMENT:long_name = "Comment applying to this parameter calibration" ;
		SCIENTIFIC_CALIB_COMMENT:_FillValue = " " ;
	char SCIENTIFIC_CALIB_DATE(N_PROF, N_CALIB, N_PARAM, DATE_TIME) ;
		SCIENTIFIC_CALIB_DATE:long_name = "Date of calibration" ;
		SCIENTIFIC_CALIB_DATE:conventions = "YYYYMMDDHHMISS" ;
		SCIENTIFIC_CALIB_DATE:_FillValue = " " ;
	char HISTORY_INSTITUTION(N_HISTORY, N_PROF, STRING4) ;
		HISTORY_INSTITUTION:long_name = "Institution which performed action" ;
		HISTORY_INSTITUTION:conventions = "Argo reference table 4" ;
		HISTORY_INSTITUTION:_FillValue = " " ;
	char HISTORY_STEP(N_HISTORY, N_PROF, STRING4) ;
		HISTORY_STEP:long_name = "Step in data processing" ;
		HISTORY_STEP:conventions = "Argo reference table 12" ;
		HISTORY_STEP:_FillValue = " " ;
	char HISTORY_SOFTWARE(N_HISTORY, N_PROF, STRING4) ;
		HISTORY_SOFTWARE:long_name = "Name of software which performed action" ;
		HISTORY_SOFTWARE:conventions = "Institution dependent" ;
		HISTORY_SOFTWARE:_FillValue = " " ;
	char HISTORY_SOFTWARE_RELEASE(N_HISTORY, N_PROF, STRING4) ;
		HISTORY_SOFTWARE_RELEASE:long_name = "Version/release of software which performed action" ;
		HISTORY_SOFTWARE_RELEASE:conventions = "Institution dependent" ;
		HISTORY_SOFTWARE_RELEASE:_FillValue = " " ;
	char HISTORY_REFERENCE(N_HISTORY, N_PROF, STRING64) ;
		HISTORY_REFERENCE:long_name = "Reference of database" ;
		HISTORY_REFERENCE:conventions = "Institution dependent" ;
		HISTORY_REFERENCE:_FillValue = " " ;
	char HISTORY_DATE(N_HISTORY, N_PROF, DATE_TIME) ;
		HISTORY_DATE:long_name = "Date the history record was created" ;
		HISTORY_DATE:conventions = "YYYYMMDDHHMISS" ;
		HISTORY_DATE:_FillValue = " " ;
	char HISTORY_ACTION(N_HISTORY, N_PROF, STRING4) ;
		HISTORY_ACTION:long_name = "Action performed on data" ;
		HISTORY_ACTION:conventions = "Argo reference table 7" ;
		HISTORY_ACTION:_FillValue = " " ;
	char HISTORY_PARAMETER(N_HISTORY, N_PROF, STRING64) ;
		HISTORY_PARAMETER:long_name = "Station parameter action is performed on" ;
		HISTORY_PARAMETER:conventions = "Argo reference table 3" ;
		HISTORY_PARAMETER:_FillValue = " " ;
	float HISTORY_START_PRES(N_HISTORY, N_PROF) ;
		HISTORY_START_PRES:long_name = "Start pressure action applied on" ;
		HISTORY_START_PRES:units = "decibar" ;
		HISTORY_START_PRES:_FillValue = 99999.f ;
	float HISTORY_STOP_PRES(N_HISTORY, N_PROF) ;
		HISTORY_STOP_PRES:long_name = "Stop pressure action applied on" ;
		HISTORY_STOP_PRES:units = "decibar" ;
		HISTORY_STOP_PRES:_FillValue = 99999.f ;
	float HISTORY_PREVIOUS_VALUE(N_HISTORY, N_PROF) ;
		HISTORY_PREVIOUS_VALUE:long_name = "Parameter/Flag previous value before action" ;
		HISTORY_PREVIOUS_VALUE:_FillValue = 99999.f ;
	char HISTORY_QCTEST(N_HISTORY, N_PROF, STRING16) ;
		HISTORY_QCTEST:long_name = "Documentation of tests performed, tests failed (in hex form)" ;
		HISTORY_QCTEST:conventions = "Write tests performed when ACTION=QCP$; tests failed when ACTION=QCF$" ;
		HISTORY_QCTEST:_FillValue = " " ;

// global attributes:
		:title = "Argo float vertical profile" ;
		:institution = "AOML" ;
		:source = "Argo float" ;
		:history = "2012-05-20 AOML 2.2 creation; 2015-05-29T19:36:21Z UW 3.1 conversion" ;
		:references = "http://www.argodatamgt.org/Documentation" ;
		:comment = "free text" ;
		:user_manual_version = "3.1" ;
		:Conventions = "Argo-3.1 CF-1.6" ;
		:featureType = "trajectoryProfile" ;
data:

 DATA_TYPE = "B-Argo profile                  " ;

 FORMAT_VERSION = "3.1 " ;

 HANDBOOK_VERSION = "1.2 " ;

 REFERENCE_DATE_TIME = "19500101000000" ;

 PLATFORM_NUMBER =
  "1900722 " ;

 PROJECT_NAME =
  "US ARGO PROJECT                                                 " ;

 PI_NAME =
  "STEPHEN RISER                                                   " ;

 STATION_PARAMETERS =
  "PRES                                                            ",
  "TEMP_DOXY                                                       ",
  "BPHASE_DOXY                                                     ",
  "DOXY                                                            " ;

 CYCLE_NUMBER = 2 ;

 DIRECTION = "A" ;

 DATA_CENTRE =
  "AO" ;

 DATE_CREATION = "20120520122653" ;

 DATE_UPDATE = "20150529123621" ;

 DC_REFERENCE =
  "1726_17964_002                  " ;

 DATA_STATE_INDICATOR =
  "2B  " ;

//********* reset P_D_M to make DATA_MODE inconsistent ***********
 DATA_MODE = "R" ;

 PARAMETER_DATA_MODE =
  "RRDR" ;

 PLATFORM_TYPE =
  "APEX                            " ;

 FLOAT_SERIAL_NO =
  "2596                            " ;

 FIRMWARE_VERSION =
  "012606                          " ;

 WMO_INST_TYPE =
  "846 " ;

 JULD = 20758.2808217439 ;

 JULD_QC = "1" ;

 JULD_LOCATION = 20758.3432986438 ;

 LATITUDE = -40.39 ;

 LONGITUDE = 73.528 ;

 POSITION_QC = "1" ;

 POSITIONING_SYSTEM =
  "ARGOS   " ;

 VERTICAL_SAMPLING_SCHEME =
  "Primary sampling: discrete []                                                                                                                                                                                                                                   " ;

 CONFIG_MISSION_NUMBER = 1 ;

 PROFILE_TEMP_DOXY_QC = " " ;

 PROFILE_BPHASE_DOXY_QC = " " ;

 PROFILE_DOXY_QC = " " ;

 PRES =
      6.5,    10.3,    20.1,    30.5,    39.7,    50.4,    60.4,    70.5, 
       80.4,    90.1,   100.0,   110.0,   120.4,   130.2,   140.4,   150.5, 
      159.8,   169.7,   180.3,   190.1,   200.2,   210.2,   220.3,   229.2, 
      240.4,   250.4,   259.5,   269.8,   279.9,   290.1,   299.6,   309.6, 
      319.7,   329.9,   339.5,   349.8,   360.2,   380.6,   400.0,   450.0, 
      500.3,   550.1,   600.4,   650.3,   700.1,   749.6,   800.3,   850.3, 
      900.1,   950.3,  1000.4,  1050.0,  1100.2,  1150.4,  1200.0,  1249.8, 
     1298.4,  1350.5,  1400.2,  1450.0,  1499.9,  1549.8,  1600.2,  1649.8, 
     1700.4,  1750.0,  1800.5,  1850.1,  1899.5,  1949.5,  1999.8 ;

 TEMP_DOXY =
     12.940,    12.940,    12.800,    12.750,    12.720,    12.710, 
       12.700,    12.680,    12.640,    12.590,    12.570,    12.550, 
       12.530,    12.510,    12.490,    12.440,    12.440,    12.430, 
       12.410,    12.360,    12.320,    12.310,    12.240,    12.170, 
       12.110,    12.070,    12.050,    12.020,    11.960,    11.940, 
       11.860,    11.760,    11.710,    11.610,    11.510,    11.380, 
       11.280,    10.900,    11.020,    10.360,    10.200,     9.750, 
        9.210,     8.740,     8.050,     7.400,     6.790,     6.120, 
        5.510,     5.140,     4.730,     4.400,     4.130,     3.840, 
        3.620,     3.520,     3.410,     3.290,     3.180,     3.080, 
        3.000,     2.910,     2.860,     2.780,     2.720,     2.670, 
        2.620,     2.590,     2.570,     2.540,     2.490 ;

 TEMP_DOXY_QC =
  "00000000000000000000000000000000000000000000000000000000000000000000000" ;

//****** add an adjusted value to a "R" variable *****
 TEMP_DOXY_ADJUSTED =
    12.940, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TEMP_DOXY_ADJUSTED_QC =
  "                                                                       " ;

 TEMP_DOXY_ADJUSTED_ERROR =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 BPHASE_DOXY =
     31.52,    31.52,    31.61,    31.66,    31.71,    31.79,    31.87, 
       31.92,    32.00,    32.12,    32.19,    32.21,    32.25,    32.28, 
       32.34,    32.45,    32.52,    32.55,    32.57,    32.62,    32.65, 
       32.73,    32.87,    32.95,    33.02,    33.07,    33.14,    33.12, 
       33.17,    33.38,    33.45,    33.46,    33.43,    33.49,    33.69, 
       33.62,    33.51,    33.43,    33.95,    34.91,    35.58,    36.18, 
       36.82,    37.38,    38.05,    38.35,    38.71,    38.61,    38.91, 
       39.30,    39.54,    39.88,    40.31,    40.83,    41.42,    41.71, 
       42.11,    42.51,    42.78,    43.06,    43.29,    43.46,    43.55, 
       43.62,    43.65,    43.65,    43.60,    43.57,    43.54,    43.46, 
       43.38 ;

 BPHASE_DOXY_QC =
  "00000000000000000000000000000000000000000000000000000000000000000000000" ;

 BPHASE_DOXY_ADJUSTED =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 BPHASE_DOXY_ADJUSTED_QC =
  "                                                                       " ;

 BPHASE_DOXY_ADJUSTED_ERROR =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 DOXY =
    231.635,   231.663,   231.275,   230.873,   230.289,   229.008, 
      227.727,   227.076,   226.064,   224.428,   223.425,   223.310, 
      222.850,   222.564,   221.763,   220.357,   219.215,   218.853, 
      218.753,   218.390,   218.294,   217.087,   215.382,   214.699, 
      214.108,   213.679,   212.748,   213.393,   213.137,   209.920, 
      209.503,   210.235,   211.206,   211.127,   208.761,   211.050, 
      213.765,   218.510,   209.043,   199.645,   191.159,   186.227, 
      181.586,   177.686,   174.020,   174.977,   174.899,   181.368, 
      182.132,   179.861,   179.946,   178.107,   174.690,   170.332, 
      164.740,   162.130,   158.316,   154.657,   152.476,   150.147, 
      148.273,   147.138,   146.657,   146.560,   146.795,   147.292, 
      148.351,   149.074,   149.742,   151.036,   152.461 ;

 DOXY_QC =
  "00000000000000000000000000000000000000000000000000000000000000000000000" ;

 DOXY_ADJUSTED =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 DOXY_ADJUSTED_QC =
  "                                                                       " ;

 DOXY_ADJUSTED_ERROR =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARAMETER =
  "PRES                                                            ",
  "TEMP_DOXY                                                       ",
  "BPHASE_DOXY                                                     ",
  "DOXY                                                            " ;

 SCIENTIFIC_CALIB_EQUATION =
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            " ;

 SCIENTIFIC_CALIB_COEFFICIENT =
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            " ;

 SCIENTIFIC_CALIB_COMMENT =
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            ",
  "none                                                                                                                                                                                                                                                            " ;

 SCIENTIFIC_CALIB_DATE =
  "              ",
  "              ",
  "              ",
  "              " ;

 HISTORY_INSTITUTION =
  "AO  " ;

 HISTORY_STEP =
  "ARFM" ;

 HISTORY_SOFTWARE =
  "    " ;

 HISTORY_SOFTWARE_RELEASE =
  "    " ;

 HISTORY_REFERENCE =
  "                                                                " ;

 HISTORY_DATE =
  "20120520122653" ;

 HISTORY_ACTION =
  "    " ;

 HISTORY_PARAMETER =
  "                                                                " ;

 HISTORY_START_PRES =
  _ ;

 HISTORY_STOP_PRES =
  _ ;

 HISTORY_PREVIOUS_VALUE =
  _ ;

 HISTORY_QCTEST =
  "                " ;
}
