netcdf argo-trajectory-v2.1-spec {

//@ DATA_TYPE = "Argo trajectory"
//@ FORMAT_VERSION   = "2.2"
//@ HANDBOOK_VERSION = "1.2"
//@ REFERENCE_DATE_TIME = "19500101000000"
//@ $Revision: 656 $
//@ $Date: 2017-04-24 16:47:02 +0000 (Mon, 24 Apr 2017) $

dimensions:
	DATE_TIME = 14;
	STRING256 = 256;
	STRING64 = 64;
	STRING32 = 32;
	STRING16 = 16;
	STRING8 = 8;
	STRING4 = 4;
	STRING2 = 2;

	N_PARAM = _unspecified_;
	N_CYCLE = _unspecified_;
	N_HISTORY = _unspecified_;
	N_HISTORY2 = _unspecified_;
	N_MEASUREMENT = UNLIMITED;

variables:
	char DATA_TYPE(STRING16);
		DATA_TYPE:comment = "Data type";
		DATA_TYPE:_FillValue = " ";
	char FORMAT_VERSION(STRING4);
		FORMAT_VERSION:comment = "File format version";
		FORMAT_VERSION:_FillValue = " ";
	char HANDBOOK_VERSION(STRING4);
		HANDBOOK_VERSION:comment = "Data handbook version";
		HANDBOOK_VERSION:_FillValue = " ";
	char REFERENCE_DATE_TIME(DATE_TIME);
		REFERENCE_DATE_TIME:comment = "Date of reference for Julian days";
		REFERENCE_DATE_TIME:conventions = "YYYYMMDDHHMISS";
		REFERENCE_DATE_TIME:_FillValue = " ";
	char PLATFORM_NUMBER(STRING8);
		PLATFORM_NUMBER:long_name = "Float unique identifier";
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII";
		PLATFORM_NUMBER:_FillValue = " ";
	char PROJECT_NAME(STRING64);
		PROJECT_NAME:comment = "Name of the project";
		PROJECT_NAME:_FillValue = " ";
	char PI_NAME (STRING64);
		PI_NAME:comment = "Name of the principal investigator";
		PI_NAME:_FillValue = " ";
	char TRAJECTORY_PARAMETERS(N_PARAM, STRING16);
		TRAJECTORY_PARAMETERS:long_name = "List of available parameters for the station";
		TRAJECTORY_PARAMETERS:conventions = "Argo reference table 3";
		TRAJECTORY_PARAMETERS:_FillValue = " ";
	char DATA_CENTRE(STRING2);
		DATA_CENTRE:long_name = "Data centre in charge of float data processing";
		DATA_CENTRE:conventions = "Argo reference table 4";
		DATA_CENTRE:_FillValue = " ";
	char DATE_CREATION(DATE_TIME);
		DATE_CREATION:comment = "Date of file creation";
		DATE_CREATION:conventions = "YYYYMMDDHHMISS";
		DATE_CREATION:_FillValue = " ";
	char DATE_UPDATE(DATE_TIME);
		DATE_UPDATE:long_name = "Date of update of this file";
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS";
		DATE_UPDATE:_FillValue = " ";
	char DATA_STATE_INDICATOR(STRING4);
		DATA_STATE_INDICATOR:long_name = "Degree of processing the data have passed through";
		DATA_STATE_INDICATOR:conventions = "Argo reference table 6";
		DATA_STATE_INDICATOR:_FillValue = " ";
	char INST_REFERENCE(STRING64);
		INST_REFERENCE:long_name = "Instrument type";
		INST_REFERENCE:conventions = "Brand, type, serial number";
		INST_REFERENCE:_FillValue = " ";
	char WMO_INST_TYPE(STRING4);
		WMO_INST_TYPE:long_name = "Coded instrument type";
		WMO_INST_TYPE:conventions = "Argo reference table 8";
		WMO_INST_TYPE:_FillValue = " ";
	char POSITIONING_SYSTEM(STRING8);
		POSITIONING_SYSTEM:long_name = "Positioning system";
		POSITIONING_SYSTEM:_FillValue = " ";
	char DATA_MODE(N_MEASUREMENT);
		DATA_MODE:long_name = "Delayed mode or real time data";
		DATA_MODE:conventions = "R : real time; D : delayed mode; A : real time with adjustment";
		DATA_MODE:_FillValue = " ";
	char DC_REFERENCE(N_MEASUREMENT, STRING32);
		DC_REFERENCE:long_name = "Location unique identifier in data centre";
		DC_REFERENCE:conventions = "Data centre convention";
		DC_REFERENCE:_FillValue = " ";
	double JULD(N_MEASUREMENT);
		JULD:long_name = "Julian day (UTC) of each measurement relative to REFERENCE_DATE_TIME";
		JULD:units = "days since 1950-01-01 00:00:00 UTC";
		JULD:conventions = "Relative julian days with decimal part (as parts of the day)";
		JULD:_FillValue = 999999.;
	char JULD_QC(N_MEASUREMENT);
		JULD_QC:long_name = "Quality on date and time";
		JULD_QC:conventions = "Argo reference table 2";
		JULD_QC:_FillValue = " ";
	double LATITUDE(N_MEASUREMENT);
		LATITUDE:long_name = "Latitude of each location";
		LATITUDE:units = "degree_north";
		LATITUDE:_FillValue = 99999.;
		LATITUDE:valid_min = -90.;
		LATITUDE:valid_max = 90.;
	double LONGITUDE(N_MEASUREMENT);
		LONGITUDE:long_name = "Longitude of each location";
		LONGITUDE:units = "degree_east";
		LONGITUDE:_FillValue = 99999.;
		LONGITUDE:valid_min = -180.;
		LONGITUDE:valid_max = 180.;
	char POSITION_ACCURACY(N_MEASUREMENT);
		POSITION_ACCURACY:long_name = "Estimated accuracy in latitude and longitude";
		POSITION_ACCURACY:conventions = "Argo reference table 5";
		POSITION_ACCURACY:_FillValue = " ";
	char POSITION_QC(N_MEASUREMENT);
		POSITION_QC:long_name = "Quality on position";
		POSITION_QC:conventions = "Argo reference table 2";
		POSITION_QC:_FillValue = " ";
	int CYCLE_NUMBER(N_MEASUREMENT);
		CYCLE_NUMBER:long_name = "Float cycle number of the measurement";
		CYCLE_NUMBER:conventions = "0..N, 0 : launch cycle, 1 : first complete cycle";
		CYCLE_NUMBER:_FillValue = 99999;

// Template (<X> indicates values from Table 3):
// Inserted based on argo-params-spec-v2.2
//	float <PARAM>(N_MEASUREMENT);
//		<PARAM>:long_name = "<X>";
//		<PARAM>:_FillValue = <X>;
//		<PARAM>:units = "<X>";
//		<PARAM>:valid_min = <X>;
//		<PARAM>:valid_max = <X>;
//		<PARAM>:comment = "<X>";
//		<PARAM>:C_format = "<X>";
//		<PARAM>:FORTRAN_format = "<X>";
//		<PARAM>:resolution = <X>;
//	char <PARAM>_QC(N_MEASUREMENT);
//		<PARAM>_QC:long_name = "quality flag";
//		<PARAM>_QC:conventions = "Argo reference table 2";
//		<PARAM>_QC:_FillValue = " ";
//	float <PARAM>_ADJUSTED(N_MEASUREMENT);
//		<PARAM>_ADJUSTED:long_name = "<X>";
//		<PARAM>_ADJUSTED:_FillValue = <X>;
//		<PARAM>_ADJUSTED:units = "<X>";
//		<PARAM>_ADJUSTED:valid_min = <X>;
//		<PARAM>_ADJUSTED:valid_max = <X>;
//		<PARAM>_ADJUSTED:comment = "<X>";
//		<PARAM>_ADJUSTED:C_format = "<X>";
//		<PARAM>_ADJUSTED:FORTRAN_format = "<X>";
//		<PARAM>_ADJUSTED:resolution= <X>;
//	char <PARAM>_ADJUSTED_QC(N_MEASUREMENT);
//		<PARAM>_ADJUSTED_QC:long_name = "quality flag";
//		<PARAM>_ADJUSTED_QC:conventions = "Argo reference table 2";
//		<PARAM>_ADJUSTED_QC:_FillValue = " ";
//	float <PARAM>_ADJUSTED_ERROR(N_MEASUREMENT);
//		<PARAM>_ADJUSTED_ERROR:long_name = "<X>";
//		<PARAM>_ADJUSTED_ERROR:_FillValue = <X>;
//		<PARAM>_ADJUSTED_ERROR:units = "<X>";
//		<PARAM>_ADJUSTED_ERROR:comment = "Contains the error on the adjusted values as determined by the delayed mode QC process.";
//		<PARAM>_ADJUSTED_ERROR:C_format = "<X>";
//		<PARAM>_ADJUSTED_ERROR:FORTRAN_format = "<X>";
//		<PARAM>_ADJUSTED_ERROR:resolution = <X>;

	double JULD_ASCENT_START(N_CYCLE);
		JULD_ASCENT_START:long_name = "Start date of the ascending profile";
		JULD_ASCENT_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_ASCENT_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_ASCENT_START:_FillValue = 999999.;
	char JULD_ASCENT_START_STATUS(N_CYCLE);
		JULD_ASCENT_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_ASCENT_START_STATUS:_FillValue = " ";
	double JULD_ASCENT_END(N_CYCLE);
		JULD_ASCENT_END:long_name = "End date of the ascending profile";
		JULD_ASCENT_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_ASCENT_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_ASCENT_END:_FillValue = 999999.;
	char JULD_ASCENT_END_STATUS(N_CYCLE);
		JULD_ASCENT_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_ASCENT_END_STATUS:_FillValue = " ";
	double JULD_DESCENT_START(N_CYCLE);
		JULD_DESCENT_START:long_name = "Descent start date of the cycle";
		JULD_DESCENT_START:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DESCENT_START:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DESCENT_START:_FillValue = 999999.;
	char JULD_DESCENT_START_STATUS(N_CYCLE);
		JULD_DESCENT_START_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DESCENT_START_STATUS:_FillValue = " ";
	double JULD_DESCENT_END(N_CYCLE);
		JULD_DESCENT_END:long_name = "Descent end date of the cycle";
		JULD_DESCENT_END:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_DESCENT_END:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_DESCENT_END:_FillValue = 999999.;
	char JULD_DESCENT_END_STATUS(N_CYCLE);
		JULD_DESCENT_END_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_DESCENT_END_STATUS:_FillValue = " ";
	double JULD_START_TRANSMISSION(N_CYCLE);
		JULD_START_TRANSMISSION:long_name = "Start date of transmission";
		JULD_START_TRANSMISSION:units = "days since 1950-01-01 00:00:00 UTC";
		JULD_START_TRANSMISSION:conventions = "Relative julian days with decimal part (as part of day)";
		JULD_START_TRANSMISSION:_FillValue = 999999.;
	char JULD_START_TRANSMISSION_STATUS(N_CYCLE);
		JULD_START_TRANSMISSION_STATUS:conventions = "0 : Nominal, 1 : Estimated, 2 : Transmitted";
		JULD_START_TRANSMISSION_STATUS:_FillValue = " ";
	char GROUNDED(N_CYCLE);
		GROUNDED:long_name = "Did the profiler touch the ground for that cycle";
		GROUNDED:conventions = "Y,N,U";
		GROUNDED:_FillValue = " ";

	char HISTORY_INSTITUTION (N_HISTORY, STRING4);
		HISTORY_INSTITUTION:long_name = "Institution which performed action";
		HISTORY_INSTITUTION:conventions = "Argo reference table 4";
		HISTORY_INSTITUTION:_FillValue = " ";
	char HISTORY_STEP(N_HISTORY, STRING4);
		HISTORY_STEP:long_name = "Step in data processing";
		HISTORY_STEP:conventions = "Argo reference table 12";
		HISTORY_STEP:_FillValue = " ";
	char HISTORY_SOFTWARE(N_HISTORY, STRING4);
		HISTORY_SOFTWARE:long_name = "Name of software which performed action";
		HISTORY_SOFTWARE:conventions = "Institution dependent";
		HISTORY_SOFTWARE:_FillValue = " ";
	char HISTORY_SOFTWARE_RELEASE(N_HISTORY, STRING4);
		HISTORY_SOFTWARE_RELEASE:long_name = "Version/release of software which performed action";
		HISTORY_SOFTWARE_RELEASE:conventions = "Institution dependent";
		HISTORY_SOFTWARE_RELEASE:_FillValue = " ";
	char HISTORY_REFERENCE(N_HISTORY, STRING64);
		HISTORY_REFERENCE:long_name = "Reference of database";
		HISTORY_REFERENCE:conventions = "Institution dependent";
		HISTORY_REFERENCE:_FillValue = " ";
	char HISTORY_DATE(N_HISTORY, DATE_TIME);
		HISTORY_DATE:long_name = "Date the history record was created";
		HISTORY_DATE:conventions = "YYYYMMDDHHMISS";
		HISTORY_DATE:_FillValue = " ";
	char HISTORY_ACTION(N_HISTORY, STRING4);
		HISTORY_ACTION:long_name = "Action performed on data";
		HISTORY_ACTION:conventions = "Argo reference table 7";
		HISTORY_ACTION:_FillValue = " ";
	char HISTORY_PARAMETER(N_HISTORY, STRING16);
		HISTORY_PARAMETER:long_name = "Station parameter action is performed on";
		HISTORY_PARAMETER:conventions = "Argo reference table 3";
		HISTORY_PARAMETER:_FillValue = " ";
	float HISTORY_PREVIOUS_VALUE(N_HISTORY, N_HISTORY2);
		HISTORY_PREVIOUS_VALUE:long_name = "Parameter/Flag previous value before action";
		HISTORY_PREVIOUS_VALUE:_FillValue = 99999.f;
        char HISTORY_INDEX_DIMENSION(N_HISTORY);
	int HISTORY_START_INDEX(N_HISTORY);
		HISTORY_START_INDEX:long_name = "Start index action applied on";
		HISTORY_START_INDEX:_FillValue = 99999;
	int HISTORY_STOP_INDEX(N_HISTORY);
		HISTORY_STOP_INDEX:long_name = "Stop index action applied on";
		HISTORY_STOP_INDEX:_FillValue = 99999;
	char HISTORY_QCTEST(N_HISTORY, N_HISTORY2, STRING16);
		HISTORY_QCTEST:long_name = "Documentation of tests performed, tests failed (in hex form)";
		HISTORY_QCTEST:conventions = "Write tests performed when ACTION=QCP$; tests failed when ACTION=QCF$";
		HISTORY_QCTEST:_FillValue = " ";
}
