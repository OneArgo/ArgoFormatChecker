netcdf argo-technical-v3.0-spec {

//@ DATA_TYPE = "Argo technical"
//@ FORMAT_VERSION   = "3.0"
//@ HANDBOOK_VERSION = "3.0"
//@ $Revision: 656 $
//@ $Date: 2017-04-24 16:47:02 +0000 (Mon, 24 Apr 2017) $

dimensions:

	DATE_TIME = 14;
	STRING128 = 128;
	STRING32 = 32;
	STRING8 = 8;
	STRING4 = 4;
	STRING2 = 2;
	N_TECH_PARAM = UNLIMITED;

variables:

	char PLATFORM_NUMBER(STRING8);
		PLATFORM_NUMBER:long_name = "Float unique identifier";
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII";
		PLATFORM_NUMBER:_FillValue = " ";
	char DATA_TYPE(STRING32); 
		DATA_TYPE:long_name = "Data type";
		DATA_TYPE:_FillValue = " ";
	char FORMAT_VERSION(STRING4);
		FORMAT_VERSION:long_name = "File format version";
		FORMAT_VERSION:_FillValue = " ";
	char HANDBOOK_VERSION(STRING4);
		HANDBOOK_VERSION:long_name = "Data handbook version";
		HANDBOOK_VERSION:_FillValue = " ";
	char DATA_CENTRE(STRING2);
		DATA_CENTRE:long_name = "Data centre in charge of float data processing";
		DATA_CENTRE:conventions = "Argo reference table 4";
		DATA_CENTRE:_FillValue = " ";
	char DATE_CREATION(DATE_TIME);
		DATE_CREATION:long_name = "Date of file creation";
		DATE_CREATION:conventions = "YYYYMMDDHHMISS";
		DATE_CREATION:_FillValue = " ";
	char DATE_UPDATE(DATE_TIME);
		DATE_UPDATE:long_name = "Date of update of this file";
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS";
		DATE_UPDATE:_FillValue = " ";
	char TECHNICAL_PARAMETER_NAME(N_TECH_PARAM, STRING128);
		TECHNICAL_PARAMETER_NAME:long_name = "Name of technical parameter";
		TECHNICAL_PARAMETER_NAME:_FillValue = " ";
	char TECHNICAL_PARAMETER_VALUE(N_TECH_PARAM, STRING128);
		TECHNICAL_PARAMETER_VALUE:long_name = "Value of technical parameter";
		TECHNICAL_PARAMETER_VALUE:_FillValue = " ";
	int CYCLE_NUMBER(N_TECH_PARAM);
		CYCLE_NUMBER:long_name = "Float cycle number";
		CYCLE_NUMBER:conventions = "0..N, 0 : launch cycle (if exists), 1 : first complete cycle";
		CYCLE_NUMBER:_FillValue = 99999;



}
