netcdf argo-metadata-v2.1-spec {

//@ DATA_TYPE = "Argo meta-data"
//@ FORMAT_VERSION   = "2.2"
//@ HANDBOOK_VERSION = "1.2"
//@ $Revision: 656 $
//@ $Date: 2017-04-24 16:47:02 +0000 (Mon, 24 Apr 2017) $

dimensions:
	DATE_TIME = 14;
	STRING256 = 256;
	STRING64 = 64;
	STRING32 = 32;
	STRING16 = 16;
	STRING8 = 8;
	STRING4 = 4;
	STRING2 = 2;
	N_CYCLES = _unspecified_;
	N_PARAM = _unspecified_;

variables:
	char DATA_TYPE(STRING16);
		DATA_TYPE:comment = "Data type";
		DATA_TYPE:_FillValue = " ";
	char FORMAT_VERSION(STRING4);
		FORMAT_VERSION:comment = "File format version";
		FORMAT_VERSION:_FillValue = " ";
	char HANDBOOK_VERSION(STRING4);
		HANDBOOK_VERSION:comment = "Data handbook version";
		HANDBOOK_VERSION:_FillValue = " ";
	char DATE_CREATION(DATE_TIME);
		DATE_CREATION:comment = "Date of file creation";
		DATE_CREATION:conventions = "YYYYMMDDHHMISS";
		DATE_CREATION:_FillValue = " ";
	char DATE_UPDATE(DATE_TIME);
		DATE_UPDATE:long_name = "Date of update of this file";
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS";
		DATE_UPDATE:_FillValue = " ";
	char PLATFORM_NUMBER(STRING8);
		PLATFORM_NUMBER:long_name = "Float unique identifier";
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII";
		PLATFORM_NUMBER:_FillValue = " ";
	char PTT(STRING256);
		PTT:long_name = "Transmission identifier (ARGOS, ORBCOMM, etc.)";
		PTT:_FillValue = " ";
	char TRANS_SYSTEM(STRING16);
		TRANS_SYSTEM:long_name = "The telecommunications system used";
		TRANS_SYSTEM:_FillValue = " ";
	char TRANS_SYSTEM_ID(STRING32);
		TRANS_SYSTEM_ID:long_name = "The program identifier used by the transmission system";
		TRANS_SYSTEM_ID:_FillValue = " ";
	char TRANS_FREQUENCY(STRING16);
		TRANS_FREQUENCY:long_name = "The frequency of transmission from the float";
		TRANS_FREQUENCY:units = "hertz";
		TRANS_FREQUENCY:_FillValue = " ";
	float TRANS_REPETITION;
		TRANS_REPETITION:long_name = "The repetition rate of transmission from the float";
		TRANS_REPETITION:units = "second";
		TRANS_REPETITION:_FillValue = 99999.f;
	char POSITIONING_SYSTEM(STRING8);
		POSITIONING_SYSTEM:long_name = "Positioning system";
		POSITIONING_SYSTEM:_FillValue = " ";
	float CLOCK_DRIFT;
		CLOCK_DRIFT:long_name = "The rate of drift of the float clock";
		CLOCK_DRIFT:units = "decisecond/day";
		CLOCK_DRIFT:_FillValue = 99999.f;
	char PLATFORM_MODEL(STRING16);
		PLATFORM_MODEL:long_name = "Model of the float";
		PLATFORM_MODEL:_FillValue = " ";
	char PLATFORM_MAKER(STRING256);
		PLATFORM_MAKER:long_name = "The name of the manufacturer";
		PLATFORM_MAKER:_FillValue = " ";
        char INST_REFERENCE(STRING64);
		INST_REFERENCE:long_name = "Instrument type";
		INST_REFERENCE:conventions = "Brand, type, serial number";
		INST_REFERENCE:_FillValue = " ";
	char WMO_INST_TYPE(STRING4);
		WMO_INST_TYPE:long_name = "Coded instrument type";
		WMO_INST_TYPE:conventions = "Argo reference table 8";
		WMO_INST_TYPE:_FillValue = " ";
	char DIRECTION;
		DIRECTION:long_name = "Direction of the profiles";
		DIRECTION:conventions = "A: ascending profiles, B: descending and ascending profiles";
		DIRECTION:_FillValue = " ";
	char PROJECT_NAME(STRING64);
		PROJECT_NAME:long_name = "The program under which the float was deployed";
		PROJECT_NAME:_FillValue = " ";
	char DATA_CENTRE(STRING2);
		DATA_CENTRE:long_name = "Data centre in charge of float real-time processing";
		DATA_CENTRE:conventions = "Argo reference table 4";
		DATA_CENTRE:_FillValue = " ";
	char PI_NAME(STRING64);
		PI_NAME:comment = "Name of the principal investigator";
		PI_NAME:_FillValue = " ";
	char ANOMALY(STRING256);
		ANOMALY:long_name = "Describe any anomalies or problems the float may have had.";
		ANOMALY:_FillValue = " ";
	char LAUNCH_DATE(DATE_TIME);
		LAUNCH_DATE:long_name = "Date (UTC) of the deployment";
		LAUNCH_DATE:conventions = "YYYYMMDDHHMISS";
		LAUNCH_DATE:_FillValue = " ";
	double LAUNCH_LATITUDE;
		LAUNCH_LATITUDE:long_name = "Latitude of the float when deployed";
		LAUNCH_LATITUDE:units = "degrees_north";
		LAUNCH_LATITUDE:_FillValue = 99999.;
		LAUNCH_LATITUDE:valid_min = -90.;
		LAUNCH_LATITUDE:valid_max = 90.;
	double LAUNCH_LONGITUDE;
		LAUNCH_LONGITUDE:long_name = "Longitude of the float when deployed";
		LAUNCH_LONGITUDE:units = "degrees_east";
		LAUNCH_LONGITUDE:_FillValue = 99999.;
		LAUNCH_LONGITUDE:valid_min = -180.;
		LAUNCH_LONGITUDE:valid_max = 180.;
	char LAUNCH_QC;
		LAUNCH_QC:long_name = "Quality on launch date, time and location";
		LAUNCH_QC:conventions = "Argo reference table 2";
		LAUNCH_QC:_FillValue = " ";
	char START_DATE(DATE_TIME);
		START_DATE:long_name = "Date (UTC) of the first descent of the float.";
		START_DATE:conventions = "YYYYMMDDHHMISS";
		START_DATE:_FillValue = " ";
	char START_DATE_QC;
		START_DATE_QC:long_name = "Quality on start date";
		START_DATE_QC:conventions = "Argo reference table 2";
		START_DATE_QC:_FillValue = " ";
	char DEPLOY_PLATFORM(STRING32);
		DEPLOY_PLATFORM:long_name = "Identifier of the deployment platform";
		DEPLOY_PLATFORM:_FillValue = " ";
	char DEPLOY_MISSION(STRING32);
		DEPLOY_MISSION:long_name = "Identifier of the mission used to deploy the float";
		DEPLOY_MISSION:_FillValue = " ";
	char DEPLOY_AVAILABLE_PROFILE_ID(STRING256);
		DEPLOY_AVAILABLE_PROFILE_ID:long_name = "Identifier of stations used to verify the first profile";
		DEPLOY_AVAILABLE_PROFILE_ID:_FillValue = " ";
	char END_MISSION_DATE (DATE_TIME);
		END_MISSION_DATE:long_name = "Date (UTC) of the end of mission of the float";
		END_MISSION_DATE:conventions = "YYYYMMDDHHMISS";
		END_MISSION_DATE:_FillValue = " ";
	char END_MISSION_STATUS;
		END_MISSION_STATUS:long_name = "Status of the end of mission of the float";
		END_MISSION_STATUS:conventions = "T:No more transmission received, R:Retrieved";
		END_MISSION_STATUS:_FillValue = " ";
	char SENSOR(N_PARAM, STRING16);
		SENSOR:long_name = "List of sensors on the float";
		SENSOR:conventions = "Argo reference table 3";
		SENSOR:_FillValue = " ";
	char SENSOR_MAKER(N_PARAM, STRING256);
		SENSOR_MAKER:long_name = "The name of the manufacturer";
		SENSOR_MAKER:_FillValue = " ";
	char SENSOR_MODEL(N_PARAM, STRING256);
		SENSOR_MODEL:long_name = "Type of sensor";
		SENSOR_MODEL:_FillValue = " ";
	char SENSOR_SERIAL_NO(N_PARAM, STRING16);
		SENSOR_SERIAL_NO:long_name = "The serial number of the sensor";
		SENSOR_SERIAL_NO:_FillValue = " ";
	char SENSOR_UNITS(N_PARAM, STRING16);
		SENSOR_UNITS:long_name = "The units of accuracy and resolution of the sensor";
		SENSOR_UNITS:_FillValue = " ";
	float SENSOR_ACCURACY(N_PARAM);
		SENSOR_ACCURACY:long_name = "The accuracy of the sensor";
		SENSOR_ACCURACY:_FillValue = 99999.f;
	float SENSOR_RESOLUTION(N_PARAM);
		SENSOR_RESOLUTION:long_name = "The resolution of the sensor";
		SENSOR_RESOLUTION:_FillValue = 99999.f;
	char PARAMETER(N_PARAM, STRING16);
		PARAMETER:long_name = "List of parameters with calibration information";
		PARAMETER:conventions = "Argo reference table 3";
		PARAMETER:_FillValue = " ";
	char PREDEPLOYMENT_CALIB_EQUATION(N_PARAM, STRING256);
		PREDEPLOYMENT_CALIB_EQUATION:long_name = "Calibration equation for this parameter";
		PREDEPLOYMENT_CALIB_EQUATION:_FillValue = " ";
	char PREDEPLOYMENT_CALIB_COEFFICIENT(N_PARAM, STRING256);
		PREDEPLOYMENT_CALIB_COEFFICIENT:long_name = "Calibration coefficients for this equation";
		PREDEPLOYMENT_CALIB_COEFFICIENT:_FillValue = " ";
	char PREDEPLOYMENT_CALIB_COMMENT(N_PARAM, STRING256);
		PREDEPLOYMENT_CALIB_COMMENT:long_name = "Comment applying to this parameter calibration";
		PREDEPLOYMENT_CALIB_COMMENT:_FillValue = " ";

	int REPETITION_RATE(N_CYCLES);
		REPETITION_RATE:long_name = "The number of times this cycle repeats";
		REPETITION_RATE:units = "number";
		REPETITION_RATE:_FillValue = 99999;
	float CYCLE_TIME(N_CYCLES);
		CYCLE_TIME:long_name = "The total time of a cycle : descent + parking + ascent + surface";
		CYCLE_TIME:units = "decimal hour";
		CYCLE_TIME:_FillValue = 99999.f;
	float PARKING_TIME(N_CYCLES);
		PARKING_TIME:long_name = "The time spent at the parking pressure";
		PARKING_TIME:units = "decimal hour";
		PARKING_TIME:_FillValue = 99999.f;
	float DESCENDING_PROFILING_TIME(N_CYCLES);
		DESCENDING_PROFILING_TIME:long_name = "The time spent sampling the descending profile";
		DESCENDING_PROFILING_TIME:units = "decimal hour";
		DESCENDING_PROFILING_TIME:_FillValue = 99999.f;
	float ASCENDING_PROFILING_TIME(N_CYCLES);
		ASCENDING_PROFILING_TIME:long_name = "The time spent sampling the ascending profile";
		ASCENDING_PROFILING_TIME:units = "decimal hour";
		ASCENDING_PROFILING_TIME:_FillValue = 99999.f;
	float SURFACE_TIME(N_CYCLES);
		SURFACE_TIME:long_name = "The time spent at the surface.";
		SURFACE_TIME:units = "decimal hour";
		SURFACE_TIME:_FillValue = 99999.f;
	float PARKING_PRESSURE(N_CYCLES);
		PARKING_PRESSURE:long_name = "The pressure of subsurface drifts";
		PARKING_PRESSURE:units = "decibar";
		PARKING_PRESSURE:_FillValue = 99999.f;
	float DEEPEST_PRESSURE(N_CYCLES);
		DEEPEST_PRESSURE:long_name = "The deepest pressure sampled in the ascending profile";
		DEEPEST_PRESSURE:units = "decibar";
		DEEPEST_PRESSURE:_FillValue = 99999.f;
	float DEEPEST_PRESSURE_DESCENDING(N_CYCLES);
		DEEPEST_PRESSURE_DESCENDING:long_name = "The deepest pressure sampled in the descending profile";
		DEEPEST_PRESSURE_DESCENDING:units = "decibar";
		DEEPEST_PRESSURE_DESCENDING:_FillValue = 99999.f;
}
