netcdf \7900685_meta {
dimensions:
	DATE_TIME = 14 ;
	STRING2 = 2 ;
	STRING4 = 4 ;
	STRING8 = 8 ;
	STRING16 = 16 ;
	STRING32 = 32 ;
	STRING64 = 64 ;
	STRING128 = 128 ;
	STRING256 = 256 ;
	STRING1024 = 1024 ;
	N_PARAM = 1 ;
	N_SENSOR = 1 ;
	N_CONFIG_PARAM = 1 ;
	N_LAUNCH_CONFIG_PARAM = 1 ;
	N_POSITIONING_SYSTEM = 1 ;
	N_TRANS_SYSTEM = 1 ;
	N_MISSIONS = UNLIMITED ; // (4 currently)
variables:
	char DATA_TYPE(STRING16) ;
		DATA_TYPE:long_name = "Data type" ;
		DATA_TYPE:conventions = "***** bad setting for this attribute *****";
		DATA_TYPE:_FillValue = " " ;
	char FORMAT_VERSION(STRING16) ;
		FORMAT_VERSION:long_name = "File format version" ;
		FORMAT_VERSION:_FillValue = " " ;
	char HANDBOOK_VERSION(STRING4) ;
		HANDBOOK_VERSION:long_name = "Data handbook version" ;
		HANDBOOK_VERSION:_FillValue = " " ;
	char DATE_CREATION(DATE_TIME) ;
		DATE_CREATION:long_name = "Date of file creation" ;
		DATE_CREATION:conventions = "YYYYMMDDHHMISS" ;
		DATE_CREATION:comment = " " ;
		DATE_CREATION:_FillValue = " " ;
	char DATE_UPDATE(DATE_TIME) ;
		DATE_UPDATE:long_name = "Date of update of this file" ;
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS" ; 
		DATE_UPDATE:_FillValue = " " ;
	char PLATFORM_NUMBER(STRING8) ;
		PLATFORM_NUMBER:long_name = "Float unique identifier" ;
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII" ;
		PLATFORM_NUMBER:_FillValue = " " ;
	char PTT(STRING256) ;
		PTT:long_name = "Transmission identifier (ARGOS, ORBCOMM, etc.)" ;
		PTT:_FillValue = " " ;
	char TRANS_SYSTEM(N_TRANS_SYSTEM, STRING16) ;
		TRANS_SYSTEM:long_name = "Telecommunications system used" ;
		TRANS_SYSTEM:_FillValue = " " ;
	char TRANS_SYSTEM_ID(N_TRANS_SYSTEM, STRING32) ;
		TRANS_SYSTEM_ID:long_name = "Program identifier used by the transmission system" ;
		TRANS_SYSTEM_ID:_FillValue = " " ;
	char TRANS_FREQUENCY(N_TRANS_SYSTEM, STRING16) ;
		TRANS_FREQUENCY:long_name = "Frequency of transmission from the float" ;
		TRANS_FREQUENCY:units = "hertz" ;
		TRANS_FREQUENCY:_FillValue = " " ;
	char POSITIONING_SYSTEM(N_POSITIONING_SYSTEM, STRING8) ;
		POSITIONING_SYSTEM:long_name = "Positioning system" ;
		POSITIONING_SYSTEM:_FillValue = " " ;
	char PLATFORM_FAMILY(STRING256) ;
		PLATFORM_FAMILY:long_name = "Category of instrument" ;
		PLATFORM_FAMILY:conventions = "Argo reference table 22" ;
		PLATFORM_FAMILY:_FillValue = " " ;
	char PLATFORM_TYPE(STRING32) ;
		PLATFORM_TYPE:long_name = "Type of float" ;
		PLATFORM_TYPE:conventions = "Argo reference table 23" ;
		PLATFORM_TYPE:_FillValue = " " ;
	char PLATFORM_MAKER(STRING256) ;
		PLATFORM_MAKER:long_name = "Name of the manufacturer" ;
		PLATFORM_MAKER:conventions = "Argo reference table 24" ;
		PLATFORM_MAKER:_FillValue = " " ;
	char FIRMWARE_VERSION(STRING32) ;
		FIRMWARE_VERSION:long_name = "Firmware version for the float" ;
		FIRMWARE_VERSION:_FillValue = " " ;
	char MANUAL_VERSION(STRING16) ;
		MANUAL_VERSION:long_name = "Manual version for the float" ;
		MANUAL_VERSION:_FillValue = " " ;
	char FLOAT_SERIAL_NO(STRING32) ;
		FLOAT_SERIAL_NO:long_name = "Serial number of the float" ;
		FLOAT_SERIAL_NO:_FillValue = " " ;
	char STANDARD_FORMAT_ID(STRING16) ;
		STANDARD_FORMAT_ID:long_name = "Standard format number to describe the data format type for each float" ;
		STANDARD_FORMAT_ID:_FillValue = " " ;
	char DAC_FORMAT_ID(STRING16) ;
		DAC_FORMAT_ID:long_name = "Format number used by the DAC to describe the data format type for each float" ;
		DAC_FORMAT_ID:_FillValue = " " ;
	char WMO_INST_TYPE(STRING4) ;
		WMO_INST_TYPE:long_name = "Coded instrument type" ;
		WMO_INST_TYPE:conventions = "Argo reference table 8" ;
		WMO_INST_TYPE:_FillValue = " " ;
	char PROJECT_NAME(STRING64) ;
		PROJECT_NAME:long_name = "Program under which the float was deployed" ;
		PROJECT_NAME:_FillValue = " " ;
	char DATA_CENTRE(STRING2) ;
		DATA_CENTRE:long_name = "Data centre in charge of float real-time processing" ;
		DATA_CENTRE:conventions = "Argo reference table 4" ;
		DATA_CENTRE:_FillValue = " " ;
	char PI_NAME(STRING64) ;
		PI_NAME:long_name = "Name of the principal investigator" ;
		PI_NAME:_FillValue = " " ;
	char ANOMALY(STRING256) ;
		ANOMALY:long_name = "Describe any anomalies or problems the float may have had" ;
		ANOMALY:_FillValue = " " ;
	char BATTERY_TYPE(STRING64) ;
		BATTERY_TYPE:long_name = "Type of battery packs in the float" ;
		BATTERY_TYPE:_FillValue = " " ;
	char BATTERY_PACKS(STRING64) ;
		BATTERY_PACKS:long_name = "Configuration of battery packs in the float" ;
		BATTERY_PACKS:_FillValue = " " ;
	char CONTROLLER_BOARD_TYPE_PRIMARY(STRING32) ;
		CONTROLLER_BOARD_TYPE_PRIMARY:long_name = "Type of primary controller board" ;
		CONTROLLER_BOARD_TYPE_PRIMARY:_FillValue = " " ;
	char CONTROLLER_BOARD_TYPE_SECONDARY(STRING32) ;
		CONTROLLER_BOARD_TYPE_SECONDARY:long_name = "Type of secondary controller board" ;
		CONTROLLER_BOARD_TYPE_SECONDARY:_FillValue = " " ;
	char CONTROLLER_BOARD_SERIAL_NO_PRIMARY(STRING32) ;
		CONTROLLER_BOARD_SERIAL_NO_PRIMARY:long_name = "Serial number of the primary controller board" ;
		CONTROLLER_BOARD_SERIAL_NO_PRIMARY:_FillValue = " " ;
	char CONTROLLER_BOARD_SERIAL_NO_SECONDARY(STRING32) ;
		CONTROLLER_BOARD_SERIAL_NO_SECONDARY:long_name = "Serial number of the secondary controller board" ;
		CONTROLLER_BOARD_SERIAL_NO_SECONDARY:_FillValue = " " ;
	char SPECIAL_FEATURES(STRING1024) ;
		SPECIAL_FEATURES:long_name = "Extra features of the float (algorithms, compressee etc.)" ;
		SPECIAL_FEATURES:_FillValue = " " ;
	char FLOAT_OWNER(STRING64) ;
		FLOAT_OWNER:long_name = "Float owner" ;
		FLOAT_OWNER:_FillValue = " " ;
	char OPERATING_INSTITUTION(STRING64) ;
		OPERATING_INSTITUTION:long_name = "Operating institution of the float" ;
		OPERATING_INSTITUTION:_FillValue = " " ;
	char CUSTOMISATION(STRING1024) ;
		CUSTOMISATION:long_name = "Float customisation, i.e. (institution and modifications)" ;
		CUSTOMISATION:_FillValue = " " ;
	char LAUNCH_DATE(DATE_TIME) ;
		LAUNCH_DATE:long_name = "Date (UTC) of the deployment" ;
		LAUNCH_DATE:conventions = "YYYYMMDDHHMISS" ;
		LAUNCH_DATE:_FillValue = " " ;
	double LAUNCH_LATITUDE ;
		LAUNCH_LATITUDE:long_name = "Latitude of the float when deployed" ;
		LAUNCH_LATITUDE:standard_name = "latitude" ;
		LAUNCH_LATITUDE:units = "degree_north" ;
		LAUNCH_LATITUDE:_FillValue = 99999. ;
		LAUNCH_LATITUDE:valid_min = -90. ;
		LAUNCH_LATITUDE:valid_max = 90. ;
		LAUNCH_LATITUDE:axis = "Y" ;
	double LAUNCH_LONGITUDE ;
		LAUNCH_LONGITUDE:long_name = "Longitude of the float when deployed" ;
		LAUNCH_LONGITUDE:standard_name = "longitude" ;
		LAUNCH_LONGITUDE:units = "degree_east" ;
		LAUNCH_LONGITUDE:_FillValue = 99999. ;
		LAUNCH_LONGITUDE:valid_min = -180. ;
		LAUNCH_LONGITUDE:valid_max = 180. ;
		LAUNCH_LONGITUDE:axis = "X" ;
	char LAUNCH_QC ;
		LAUNCH_QC:long_name = "Quality on launch date, time and location" ;
		LAUNCH_QC:conventions = "Argo reference table 2" ;
		LAUNCH_QC:_FillValue = " " ;
	char START_DATE(DATE_TIME) ;
		START_DATE:long_name = "Date (UTC) of the first descent of the float" ;
		START_DATE:conventions = "YYYYMMDDHHMISS" ;
		START_DATE:_FillValue = " " ;
	char START_DATE_QC ;
		START_DATE_QC:long_name = "Quality on start date" ;
		START_DATE_QC:conventions = "Argo reference table 2" ;
		START_DATE_QC:_FillValue = " " ;
	char STARTUP_DATE(DATE_TIME) ;
		STARTUP_DATE:long_name = "Date (UTC) of the activation of the float" ;
		STARTUP_DATE:conventions = "YYYYMMDDHHMISS" ;
		STARTUP_DATE:_FillValue = " " ;
	char STARTUP_DATE_QC ;
		STARTUP_DATE_QC:long_name = "Quality on startup date" ;
		STARTUP_DATE_QC:conventions = "Argo reference table 2" ;
		STARTUP_DATE_QC:_FillValue = " " ;
	char DEPLOYMENT_PLATFORM(STRING32) ;
		DEPLOYMENT_PLATFORM:long_name = "Identifier of the deployment platform" ;
		DEPLOYMENT_PLATFORM:_FillValue = " " ;
	char DEPLOYMENT_CRUISE_ID(STRING32) ;
		DEPLOYMENT_CRUISE_ID:long_name = "Identification number or reference number of the cruise used to deploy the float" ;
		DEPLOYMENT_CRUISE_ID:_FillValue = " " ;
	char DEPLOYMENT_REFERENCE_STATION_ID(STRING256) ;
		DEPLOYMENT_REFERENCE_STATION_ID:long_name = "Identifier or reference number of co-located stations used to verify the first profile" ;
		DEPLOYMENT_REFERENCE_STATION_ID:_FillValue = " " ;
	char END_MISSION_DATE(DATE_TIME) ;
		END_MISSION_DATE:long_name = "Date (UTC) of the end of mission of the float" ;
		END_MISSION_DATE:conventions = "YYYYMMDDHHMISS" ;
		END_MISSION_DATE:_FillValue = " " ;
	char END_MISSION_STATUS ;
		END_MISSION_STATUS:long_name = "Status of the end of mission of the float" ;
		END_MISSION_STATUS:conventions = "T:No more transmission received, R:Retrieved" ;
		END_MISSION_STATUS:_FillValue = " " ;
	char LAUNCH_CONFIG_PARAMETER_NAME(N_LAUNCH_CONFIG_PARAM, STRING128) ;
		LAUNCH_CONFIG_PARAMETER_NAME:long_name = "Name of configuration parameter at launch" ;
		LAUNCH_CONFIG_PARAMETER_NAME:_FillValue = " " ;
	double LAUNCH_CONFIG_PARAMETER_VALUE(N_LAUNCH_CONFIG_PARAM) ;
		LAUNCH_CONFIG_PARAMETER_VALUE:long_name = "Value of configuration parameter at launch" ;
		LAUNCH_CONFIG_PARAMETER_VALUE:_FillValue = 99999. ;
	char CONFIG_PARAMETER_NAME(N_CONFIG_PARAM, STRING128) ;
		CONFIG_PARAMETER_NAME:long_name = "Name of configuration parameter" ;
		CONFIG_PARAMETER_NAME:_FillValue = " " ;
	double CONFIG_PARAMETER_VALUE(N_MISSIONS, N_CONFIG_PARAM) ;
		CONFIG_PARAMETER_VALUE:long_name = "Value of configuration parameter" ;
		CONFIG_PARAMETER_VALUE:_FillValue = 99999. ;
	int CONFIG_MISSION_NUMBER(N_MISSIONS) ;
		CONFIG_MISSION_NUMBER:long_name = "Unique number denoting the missions performed by the float" ;
		CONFIG_MISSION_NUMBER:conventions = "1...N, 1 : first complete mission" ;
		CONFIG_MISSION_NUMBER:_FillValue = 99999 ;
	char CONFIG_MISSION_COMMENT(N_MISSIONS, STRING256) ;
		CONFIG_MISSION_COMMENT:long_name = "Comment on configuration" ;
		CONFIG_MISSION_COMMENT:_FillValue = " " ;
	char SENSOR(N_SENSOR, STRING32) ;
		SENSOR:long_name = "Name of the sensor mounted on the float" ;
		SENSOR:conventions = "Argo reference table 25" ;
		SENSOR:_FillValue = " " ;
	char SENSOR_MAKER(N_SENSOR, STRING256) ;
		SENSOR_MAKER:long_name = "Name of the sensor manufacturer" ;
		SENSOR_MAKER:conventions = "Argo reference table 26" ;
		SENSOR_MAKER:_FillValue = " " ;
	char SENSOR_MODEL(N_SENSOR, STRING256) ;
		SENSOR_MODEL:long_name = "Type of sensor" ;
		SENSOR_MODEL:conventions = "Argo reference table 27" ;
		SENSOR_MODEL:_FillValue = " " ;
	char SENSOR_SERIAL_NO(N_SENSOR, STRING16) ;
		SENSOR_SERIAL_NO:long_name = "Serial number of the sensor" ;
		SENSOR_SERIAL_NO:_FillValue = " " ;
	char PARAMETER(N_PARAM, STRING64) ;
		PARAMETER:long_name = "Name of parameter computed from float measurements" ;
		PARAMETER:conventions = "Argo reference table 3" ;
		PARAMETER:_FillValue = " " ;
	char PARAMETER_SENSOR(N_PARAM, STRING128) ;
		PARAMETER_SENSOR:long_name = "Name of the sensor that measures this parameter" ;
		PARAMETER_SENSOR:conventions = "Argo reference table 25" ;
		PARAMETER_SENSOR:_FillValue = " " ;
	char PARAMETER_UNITS(N_PARAM, STRING32) ;
		PARAMETER_UNITS:long_name = "Units of accuracy and resolution of the parameter" ;
		PARAMETER_UNITS:_FillValue = " " ;
	char PARAMETER_ACCURACY(N_PARAM, STRING32) ;
		PARAMETER_ACCURACY:long_name = "Accuracy of the parameter" ;
		PARAMETER_ACCURACY:_FillValue = " " ;
	char PARAMETER_RESOLUTION(N_PARAM, STRING32) ;
		PARAMETER_RESOLUTION:long_name = "Resolution of the parameter" ;
		PARAMETER_RESOLUTION:_FillValue = " " ;
	char PREDEPLOYMENT_CALIB_EQUATION(N_PARAM, STRING1024) ;
		PREDEPLOYMENT_CALIB_EQUATION:long_name = "Calibration equation for this parameter" ;
		PREDEPLOYMENT_CALIB_EQUATION:_FillValue = " " ;
	char PREDEPLOYMENT_CALIB_COEFFICIENT(N_PARAM, STRING1024) ;
		PREDEPLOYMENT_CALIB_COEFFICIENT:long_name = "Calibration coefficients for this equation" ;
		PREDEPLOYMENT_CALIB_COEFFICIENT:_FillValue = " " ;
	char PREDEPLOYMENT_CALIB_COMMENT(N_PARAM, STRING1024) ;
		PREDEPLOYMENT_CALIB_COMMENT:long_name = "Comment applying to this parameter calibration" ;
		PREDEPLOYMENT_CALIB_COMMENT:_FillValue = " " ;

// global attributes:
		:title = "Argo float metadata file" ;
		:institution = "Scripps Institution of Oceanography" ;
		:source = "Argo float" ;
		:history = "2018-03-08T20:35:37Z creation; 2018-04-10T22:21:06Z most recent update" ;
		:references = "http://www.argodatamgt.org/Documentation" ;
		:comment = "free text" ;
		:user_manual_version = "3.10" ;
		:Conventions = "Argo-3.1 CF-1.6" ;
		:comment_on_dac_decoder_version = "Decoded by SIO: Argo SIO SOLOII V2.4" ;

data:

 DATA_TYPE = "Argo meta-data  " ;

 FORMAT_VERSION = "10.0 " ;

 HANDBOOK_VERSION = "1.2 " ;

 DATE_CREATION = "20180308203537" ;

 DATE_UPDATE = "20180410222106" ;

 PLATFORM_NUMBER = "7900685 " ;

 PTT = "n/a                                                                                                                                                                                                                                                             " ;

 TRANS_SYSTEM =
  "IRIDIUM         " ;

 TRANS_SYSTEM_ID =
  "n/a                             " ;

 TRANS_FREQUENCY =
  "n/a             " ;

 POSITIONING_SYSTEM =
  "GPS     " ;

 PLATFORM_FAMILY = "FLOAT                                                                                                                                                                                                                                                           " ;

 PLATFORM_TYPE = "SOLO_II                         " ;

 PLATFORM_MAKER = "SIO_IDG                                                                                                                                                                                                                                                         " ;

 FIRMWARE_VERSION = "V02.40; SBE602 15Aug17          " ;

 MANUAL_VERSION = "V02.40          " ;

 FLOAT_SERIAL_NO = "8637                            " ;

 STANDARD_FORMAT_ID = "202024          " ;

 DAC_FORMAT_ID = "SOLO2IR_TS36    " ;

 WMO_INST_TYPE = "853 " ;

 PROJECT_NAME = "US ARGO PROJECT                                                 " ;

 DATA_CENTRE = "AO" ;

 PI_NAME = "DEAN ROEMMICH                                                   " ;

 ANOMALY = "                                                                                                                                                                                                                                                                " ;

 BATTERY_TYPE = "Lithium                                                         " ;

 BATTERY_PACKS = "1 CPU (sn=2511); 3 PUMP (sn=17212 17208 17);                    " ;

 CONTROLLER_BOARD_TYPE_PRIMARY = "GG32 Rev:6.2                    " ;

 CONTROLLER_BOARD_TYPE_SECONDARY = "                                " ;

 CONTROLLER_BOARD_SERIAL_NO_PRIMARY = "2496                            " ;

 CONTROLLER_BOARD_SERIAL_NO_SECONDARY = "                                " ;

}
