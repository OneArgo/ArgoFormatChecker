netcdf \7900685_meta {
dimensions:
	DATE_TIME = 14 ;
	STRING2 = 2 ;
	STRING4 = 4 ;
	STRING8 = 8 ;
	STRING16 = 16 ;
	STRING32 = 32 ;
	STRING64 = 64 ;
	STRING128 = 128 ;
	STRING256 = 256 ;
	STRING1024 = 1024 ;
	N_PARAM = 3 ;
	N_SENSOR = 3 ;
	N_CONFIG_PARAM = 20 ;
	N_LAUNCH_CONFIG_PARAM = 27 ;
	N_POSITIONING_SYSTEM = 1 ;
	N_TRANS_SYSTEM = 1 ;
	N_MISSIONS = UNLIMITED ; // (4 currently)
variables:
	char DATA_TYPE(STRING16) ;
		DATA_TYPE:long_name = "Data type" ;
		DATA_TYPE:conventions = "Argo reference table 1" ;
		DATA_TYPE:_FillValue = " " ;
data:

 DATA_TYPE = "Argo meta-data  " ;

}
